library verilog;
use verilog.vl_types.all;
entity registrador1b is
    port(
        clock           : in     vl_logic;
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end registrador1b;
